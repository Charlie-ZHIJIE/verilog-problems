`timescale 1ns/1ps

module simple_adder (
    input wire clk,
    input wire [7:0] a,
    input wire [7:0] b,
    output reg [7:0] sum
);
    // TODO: Implement the adder logic
endmodule
